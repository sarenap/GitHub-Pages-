// Code your design here
`include "light_package.sv"
`include "traffic_light_controller1.sv"
