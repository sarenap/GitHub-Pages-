// Code your testbench here
// or browse Examples
`include "lab3_part1_tb.sv"
//`include "light_package.sv"